module wallace_tree_32 #(
    parameter WIDTH = 32;
) 
(
    input wire logic[WIDTH - 1:0] a,
    input wire logic[WIDTH - 1:0] b,
    output logic;WIDTH - 1:0] result,
    output logic overflow
);



endmodule