import riscv_core_p::*;

module riscv_basic_pipeline 
#(
    parameter PC_INITIAL = 0x00400000,
    parameter XLEN = 32
) (
    input wire logic clk,
    input wire logic rst,
    output logic[XLEN - 1:0] PC,
    input logic[RISCV_INSTR_LEN - 1] instruction,
    output wire logic[XLEN - 1:0] ALUResult,
    output wire logic[XLEN - 1:0] dAddress,
    output wire logic[XLEN - 1:0] dWriteData,
    output wire logic[XLEN - 1:0] dReadData,
    output wire logic MemRead,
    output wire logic MemWrite,
    output wire logic[XLEN - 1:0] WriteBackData
);

//////////////////////////////////////////////////////////////////////
// IF: Instruction Fetch
//////////////////////////////////////////////////////////////////////	



//////////////////////////////////////////////////////////////////////
// ID: Instruction Decode
//////////////////////////////////////////////////////////////////////	



//////////////////////////////////////////////////////////////////////
// EX: Execute
//////////////////////////////////////////////////////////////////////	



//////////////////////////////////////////////////////////////////////
// MEM: Memory Access
//////////////////////////////////////////////////////////////////////	


//////////////////////////////////////////////////////////////////////
// WB: Write Back
//////////////////////////////////////////////////////////////////////	


endmodule